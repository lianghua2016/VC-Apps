module top(input wire top_clk);
dut inst(top_clk);
endmodule

module dut(input wire sub_clk);
endmodule
