module dut();
endmodule

module top;
dut inst1();
dut inst2();
endmodule


